/* CSED273 lab2 experiment 2 */
/* lab2_2.v */

/* Simplifed equation by K-Map method
 * You are allowed to use keword "assign" and operator "&","|","~",
 * or just implement with gate-level-modeling (and, or, not) */
module lab2_2(
    output wire outGT, outEQ, outLT,
    input wire [1:0] inA,
    input wire [1:0] inB
    );

    CAL_GT_2 cal_gt2(outGT, inA, inB);
    CAL_EQ_2 cal_eq2(outEQ, inA, inB);
    CAL_LT_2 cal_lt2(outLT, inA, inB);

endmodule

/* Implement output about "A>B" */
module CAL_GT_2(
    output wire outGT,
    input wire [1:0] inA,
    input wire [1:0] inB
    );

    ////////////////////////
    /* Add your code here */
    // outGT�� inA�� �ֻ��� ��Ʈ�� inB�� �ֻ��� ��Ʈ���� Ŭ ��, Ȥ��
    // �ֻ��� ��Ʈ�� �����ϰ� inA�� ������ ��Ʈ�� inB�� ������ ��Ʈ���� Ŭ �� ���̴�
    assign outGT = (inA[1] & ~inB[1]) | (~inB[1] & inA[0] & ~inB[0]);
    ////////////////////////

endmodule

/* Implement output about "A=B" */
module CAL_EQ_2(
    output wire outEQ,
    input wire [1:0] inA, 
    input wire [1:0] inB
    );

    ////////////////////////
    /* Add your code here */
    // outEQ�� inA�� inB�� ��� ��Ʈ�� ��ġ�� �� ��
    // XOR ���� ����� 0�̸� �� ��Ʈ�� ���ٴ� ���� �ǹ��ϹǷ�, ���⼭�� ���� �����ڸ� ����Ѵ�
    assign outEQ = ((inA[1] ~^ inB[1]) & (inA[0] ~^ inB[0]));
    ////////////////////////

endmodule

/* Implement output about "A<B" */
module CAL_LT_2(
    output wire outLT,
    input wire [1:0] inA, 
    input wire [1:0] inB
    );

    ////////////////////////
    /* Add your code here */
    // outLT�� inA�� �ֻ��� ��Ʈ�� inB�� �ֻ��� ��Ʈ���� ���� ��, Ȥ��
    // �ֻ��� ��Ʈ�� �����ϰ� inA�� ������ ��Ʈ�� inB�� ������ ��Ʈ���� ���� �� ���Դϴ�.
    assign outLT = (~inA[1] & inB[1]) | (~inA[1] & ~inA[0] & inB[0]);
    ////////////////////////

endmodule